// GENERATE INPLACE BEGIN fileheader() =========================================
//
// GENERATE INPLACE END fileheader =============================================

// GENERATE INPLACE BEGIN beginmod() ===========================================
// GENERATE INPLACE END beginmod ===============================================

// GENERATE INPLACE BEGIN endmod() =============================================
// GENERATE INPLACE END endmod =================================================
